--Steven Miller
--11710
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity clk_gen is
    generic (
        ms_period : positive := 1000);          -- amount of ms for button to be
                                        -- pressed before creating clock pulse
    port (
        clk50MHz : in  std_logic;
        rst      : in  std_logic;
        button_n : in  std_logic;
        clk_out  : out std_logic);
end clk_gen;

architecture arch of clk_gen is
component clk_div
	generic(clk_in_freq: positive := 50000000; clk_out_freq : positive:= 1000);
	port(
		clk_in : in std_logic;
		clk_out : out std_logic;
		rst : in std_logic
	);
end component;

signal slowclk : std_logic;
begin
--modify data you feed into your divider so each count is 1 ms long
clkdiv: clk_div generic map (clk_in_freq => 50000000, clk_out_freq => 2000)
 port map(clk_in => clk50Mhz, clk_out => slowclk, rst=>rst);
process(slowclk, rst)
variable count : natural := 0;
begin
--if reset
if(rst = '1') then
	clk_out <= '0';
	count := 0;
elsif(slowclk'Event and slowclk = '1') then
	--if button held down
	if(button_n = '0') then
		--if ms_period/1000 second(s) has elapsed
		if(count = ms_period) then
			clk_out <= '1'; -- end pulse
			count := 0;
		else
			count := count +1;
			clk_out <= '0';
		end if;
	else
		clk_out <= '0';
		count := 0;
	end if;
end if;
end process;
end arch;