--Steven Miller
--11710
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.NUMERIC_STD.UNSIGNED;

entity gray2_tb is
end gray2_tb;

architecture TB of gray2_tb is

signal clk    : std_logic:='0';
signal rst : std_logic:='0';
signal output  : std_logic_vector(3 downto 0);

signal done : std_logic := '0';
begin  -- TB

  UUT : entity work.gray2
    port map 
(
      clk     => clk,
      rst     => rst,
      output  => output
);
 
clk <= not(clk) after 10 ns when done = '0' else clk;
 process

    function graycounter 
    (
      constant count      : integer
    )
      return std_logic_vector is
    begin
      case count is
	when 0 =>
		return "0000";
	when 1 =>
		return "0001";
	when 2 =>
		return "0011";
	when 3 =>
		return "0010";
	when 4 => 
		return "0110";
	when 5 =>
		return "0111";
	when 6 =>
		return "0101";
	when 7 =>
		return "0100";
	when 8 =>
		return "1100";
	when 9 =>
		return "1101";
	when 10 =>
		return "1111";
	when 11 =>
		return "1110";
	when 12 =>
		return "1010";
	when 13 =>
		return "1011";
	when 14 =>
		return "1001";
	when 15 =>
		return "1000";
	when others =>
		return "0000";
      end case;
    end graycounter;

  begin
    rst <= '1'; 
    wait for 200 ns;
    -- test count
    rst <= '0';
    wait for 200 ns;
    for i in 1 to 15 loop
	wait for 20 ns;
	assert(output = graycounter(i)) report "counter incorrect";
	wait until rising_edge(clk);
    end loop;

   --wrap back to 0 test
    wait for 10 ns;
    assert(output = graycounter(0)) report "wrap back to 0 incorrect";

   for i in 0 to 4 loop
	wait until rising_edge(clk);
    end loop;
    --reset test
    rst    <= '1';
    wait for 10 ns;
    assert(output = graycounter(0)) report "Clear failed" severity warning;
    wait for 20 ns;
    report "SIMULATION FINISHED!";
    done <= '1';

  end process;
end TB;
